-- fichier à écraser avec le fichier généré par ISE (New Source)
